module SramArbiter(
  // Application interface
  input reset,

  // W0
  input         w0_clock,
  output        w0_din_ready,
  input         w0_din_valid,
  input [53:0]  w0_din,// {mask,addr,data}

  // W1
  input         w1_clock,
  output        w1_din_ready,
  input         w1_din_valid,
  input [53:0]  w1_din,// {mask,addr,data}

  // R0
  input         r0_clock,
  output        r0_din_ready,
  input         r0_din_valid,
  input  [17:0] r0_din, // addr
  input         r0_dout_ready,
  output        r0_dout_valid,
  output [31:0] r0_dout, // data

  // R1
  input         r1_clock,
  output        r1_din_ready,
  input         r1_din_valid,
  input  [17:0] r1_din, // addr
  input         r1_dout_ready,
  output        r1_dout_valid,
  output [31:0] r1_dout, // data

  `ifdef MODELSIM // Output for testbench
  output reg [2:0] state;
  `endif

  // SRAM Interface
  input         sram_clock,
  output        sram_addr_valid, // assigned
  input         sram_ready, //TODO WHAT TO DO WITH THIS?
  output [17:0] sram_addr,
  output [31:0] sram_data_in, // assigned
  output  [3:0] sram_write_mask, // assigned
  input  [31:0] sram_data_out,
  input         sram_data_out_valid);

// Clock crossing FIFOs --------------------------------------------------------

// The SRAM_WRITE_FIFOis have been instantiated for you, but you must wire it
// correctly

localparam DOW0 = 3'b000,
           DOW1 = 3'b001,
           DOR0 = 3'b010,
           DOR1 = 3'b011,
           PAUSE = 3'b100;


reg [2:0] readshift; // potential for off by one error - might need to be 3:0
reg [2:0] CurrentState;
reg [2:0] NextState;


wire w0_valid;
wire w1_valid;

reg next2;
reg this0; // current cycle's read (only "valid" if this is a read)
reg this1;
reg this2;



wire w0_rd_en, w1_rd_en;
wire w0empty, w1empty;
wire [53:0] w0dout, w1dout;

wire r0_data_write, r1_data_write;

wire r0_data_full, r1_data_full;

wire r0_read_valid, r1_read_valid;
wire r0_addr, r1_addr;

wire r0_rd_en, r1_rd_en;




// following 3 lines handle correctly asserting w0_din_ready and w1_din_ready
wire w0_full, w1_full;
assign w0_din_ready = !w0_full;
assign w1_din_ready = !w1_full;

assign w0_rd_en = (CurrentState == DOW0);
assign w1_rd_en = (CurrentState == DOW1);

//this is fine because we don't care what's on the sram_data_in line on R0 and R1
assign sram_data_in = (CurrentState == DOW0) ? w0dout[31:0] : w1dout[31:0];
assign sram_write_mask = (CurrentState == DOW0) ? w0dout[53:50] : ((CurrentState == DOW1) ? w1dout[53:50] : 4'b0000);
assign sram_addr = (CurrentState == DOW0) ? w0dout[49:32] : ((CurrentState == DOW1) ? w1dout[49:32] : ((CurrentState == DOR0) ? r0_addr : ((CurrentState == DOR1) ? r1_addr : 0)));
assign sram_addr_valid = (CurrentState == DOW0 || CurrentState == DOW1 || CurrentState == DOR0 || CurrentState == DOR1);

SRAM_WRITE_FIFO w0_fifo(
  .rst(reset),
  .wr_clk(w0_clock),
  .din(w0_din),
  .wr_en(w0_din_valid),
  .full(w0_full),

  .rd_clk(sram_clock), //sram_clock is our "internal clock"
  .rd_en(w0_rd_en),
  .valid(w0_valid),
  .dout(w0dout),
  .empty()); // unused?

SRAM_WRITE_FIFO w1_fifo(
  .rst(reset),
  .wr_clk(w1_clock),
  .din(w1_din),
  .wr_en(w1_din_valid),
  .full(w1_full),

  .rd_clk(sram_clock), //sram_clock is our "internal clock"
  .rd_en(w1_rd_en),
  .valid(w1_valid),
  .dout(w1dout),
  .empty()); // unused?


// Instantiate the Read FIFOs here
assign r0_data_write = sram_data_out_valid & (!this0);
assign r1_data_write = sram_data_out_valid & this0;


SRAM_DATA_FIFO r0_data_fifo(
  .rst(reset),
  .wr_clk(sram_clock),
  .din(sram_data_out),
  .wr_en(r0_data_write),
  .full(),

  .rd_clk(r0_clock),
  .rd_en(r0_dout_ready),
  .valid(r0_dout_valid),
  .dout(r0_dout),
  .empty(),
  .prog_full());


SRAM_DATA_FIFO r1_data_fifo(
  .rst(reset),
  .wr_clk(sram_clock),
  .din(sram_data_out),
  .wr_en(r1_data_write),
  .full(),

  .rd_clk(r1_clock),
  .rd_en(r1_dout_ready),
  .valid(r1_dout_valid),
  .dout(r1_dout),
  .empty(),
  .prog_full());

assign r0_din_ready = !r0_data_full; // TODO: backpressure
assign r1_din_ready = !r1_data_full; // TODO: backpressure
assign r0_rd_en = (CurrentState == DOR0);
assign r1_rd_en = (CurrentState == DOR1);

SRAM_ADDR_FIFO r0_addr_fifo(
  .rst(reset),
  .wr_clk(r0_clock),
  .din(r0_din),
  .wr_en(r0_din_valid),
  .full(r0_data_full),

  .rd_clk(sram_clock),
  .rd_en(r0_rd_en),
  .valid(r0_read_valid),
  .dout(r0_addr),
  .empty()); //unused?

SRAM_ADDR_FIFO r1_addr_fifo(
  .rst(reset),
  .wr_clk(r1_clock),
  .din(r1_din),
  .wr_en(r1_din_valid),
  .full(r1_data_full),

  .rd_clk(sram_clock),
  .rd_en(r0_rd_en),
  .valid(r1_read_valid),
  .dout(r1_addr),
  .empty()); //unused?


// Arbiter Logic ---------------------------------------------------------------

`ifdef MODELSIM // Output for testbench
always @(*)
  if (currentState == DOW0) state = 3'b00;
  else if (currentState == DOW1) state = 3'b001;
  else if (currentState == DOR0) state = 3'b010;
  else if (currentState == DOR1) state = 3'b011;
  else if (currentState == PAUSE) state = 3'b100;
  else state = 3'b111;
`endif

// need reg to keep track of whether or not a read is supposed to happen next
// cycle


always @(posedge sram_clock) begin
    if (reset) begin
        CurrentState <= PAUSE;
        this0 <= 1'b0;
        this1 <= 1'b0;
        this2 <= 1'b0;
    end
    else begin
        CurrentState <= NextState;
        this0 <= this1;
        this1 <= this2;
        this2 <= next2;
    end
end


always @(*) begin
    case(CurrentState) 
        PAUSE: begin
            if(w0_valid) NextState = DOW0;
            else if(w1_valid) NextState = DOW1;
            else if( r0_read_valid ) NextState = DOR0;
            else if( r1_read_valid ) NextState = DOR1;
            else NextState = PAUSE;
        end

        DOW0: begin
            if(w1_valid) NextState = DOW1;
            else if( r0_read_valid ) NextState = DOR0;
            else if( r1_read_valid ) NextState = DOR1;
            else if(w0_valid) NextState = DOW0;
            else NextState = PAUSE;
        end

        DOW1: begin
            if( r0_read_valid ) NextState = DOR0;
            else if( r1_read_valid ) NextState = DOR1;
            else if(w0_valid) NextState = DOW0;
            else if(w1_valid) NextState = DOW1;
            else NextState = PAUSE;
        end

        DOR0: begin
            next2 = 1'b0;
            if( r1_read_valid ) NextState = DOR1;
            else if(w0_valid) NextState = DOW0;
            else if(w1_valid) NextState = DOW1;
            else if( r0_read_valid ) NextState = DOR0;
            else NextState = PAUSE;
        end

        DOR1: begin
            next2 = 1'b1;
            if(w0_valid) NextState = DOW0;
            else if(w1_valid) NextState = DOW1;
            else if( r0_read_valid ) NextState = DOR0;
            else if( r1_read_valid ) NextState = DOR1;
            else NextState = PAUSE;
        end

    endcase
end

// Put your round-robin arbitration logic here

endmodule
